LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MY_CIRCUIT2 IS
	PORT (S: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
	      D: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
              Y: OUT STD_LOGIC);
END MY_CIRCUIT2;

ARCHITECTURE MY_CIRCUIT_ARCH2 OF MY_CIRCUIT2 IS
BEGIN
	Y <= (D(0) AND NOT(S(1)) AND NOT(S(0))) OR (D(1) AND NOT(S(1)) AND S(0)) OR (D(2) AND S(1) AND NOT(S(0))) OR (D(3) AND S(1) AND S(0));
END MY_CIRCUIT_ARCH2;