LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SOMADOR_PALAVRAS_4BITS IS
    PORT(A : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
         B : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
         S : OUT STD_LOGIC_VECTOR(4 DOWNTO 0));
END ENTITY SOMADOR_PALAVRAS_4BITS;

ARCHITECTURE SOMADOR_PALAVRAS_4BITS_ARCH OF SOMADOR_PALAVRAS_4BITS IS

    COMPONENT SOMADOR_COMPLETO IS
        PORT(A, B, CIN : IN  STD_LOGIC;
             S, COUT   : OUT STD_LOGIC);
    END COMPONENT;

    SIGNAL COUT0, COUT1, COUT2 : STD_LOGIC;

BEGIN

    SOMADOR0: SOMADOR_COMPLETO
        PORT MAP(A => A(0), B => B(0), CIN => '0',   S => S(0), COUT => COUT0);

    SOMADOR1: SOMADOR_COMPLETO
        PORT MAP(A => A(1), B => B(1), CIN => COUT0, S => S(1), COUT => COUT1);

    SOMADOR2: SOMADOR_COMPLETO
        PORT MAP(A => A(2), B => B(2), CIN => COUT1, S => S(2), COUT => COUT2);

    SOMADOR3: SOMADOR_COMPLETO
        PORT MAP(A => A(3), B => B(3), CIN => COUT2, S => S(3), COUT => S(4));

END ARCHITECTURE SOMADOR_PALAVRAS_4BITS_ARCH;

