LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY TB_SOMADORPALAVRAS IS
END ENTITY;

ARCHITECTURE behavior OF TB_SOMADORPALAVRAS IS
    SIGNAL A_TB, B_TB : STD_LOGIC_VECTOR(3 DOWNTO 0);
    SIGNAL S_TB       : STD_LOGIC_VECTOR(4 DOWNTO 0);
BEGIN
    UUT: ENTITY WORK.SOMADORPALAVRAS
        PORT MAP(
            A => A_TB,
            B => B_TB,
            S => S_TB
        );

    PROCESS
    BEGIN
        A_TB <= "0000"; B_TB <= "0000"; WAIT FOR 10 ns;
        A_TB <= "0001"; B_TB <= "0010"; WAIT FOR 10 ns;
        A_TB <= "0111"; B_TB <= "0001"; WAIT FOR 10 ns;
        A_TB <= "1111"; B_TB <= "1111"; WAIT FOR 10 ns;

        WAIT;
    END PROCESS;
END ARCHITECTURE behavior;

