LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY GOLDENSOMADOR IS
PORT (
A,B : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
S: OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
);
END ENTITY GOLDENSOMADOR;

ARCHITECTURE GOLDENMODEL OF GOLDENSOMADOR IS
BEGIN
S <= (UNSIGNED('0' & A) + UNSIGNED('0' & B));


END GOLDENMODEL;
