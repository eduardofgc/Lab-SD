LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MY_CIRCUIT IS
	PORT (A, B, CIN: IN STD_LOGIC;
              S, COUT: OUT STD_LOGIC);
END MY_CIRCUIT;

ARCHITECTURE MY_CIRCUIT_ARCH OF MY_CIRCUIT IS
BEGIN
	S <= A XOR B XOR CIN;
        COUT <= (A AND B) OR (A AND CIN) OR (B AND CIN); 
END MY_CIRCUIT_ARCH;
