LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MY_CIRCUIT3 IS
	PORT (A: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
	      S: OUT STD_LOGIC);
END MY_CIRCUIT3;

ARCHITECTURE MY_CIRCUIT_ARCH3 OF MY_CIRCUIT3 IS
BEGIN
	S <= (A(3) AND A(2) AND NOT(A(1)) AND NOT(A(0))) OR (A(3) AND NOT(A(2)) AND NOT(A(1)) AND A(0)) OR (NOT(A(3)) AND A(2) AND NOT(A(1)) AND A(0)) OR (NOT(A(3)) AND NOT(A(2)) AND A(1) AND A(0)) OR (NOT(A(3)) AND A(2) AND A(1) AND NOT(A(0))) OR (A(3) AND A(2) AND A(1) AND A(0)) OR (A(3) AND NOT(A(2)) AND A(1) AND NOT(A(0)));
END MY_CIRCUIT_ARCH3;