LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SOMADOR IS
	PORT (A, B, CIN: IN STD_LOGIC;
              S, COUT: OUT STD_LOGIC);
END SOMADOR;

ARCHITECTURE SOMADOR_ARCH OF SOMADOR IS
BEGIN
	S <= A XOR B XOR CIN;
        COUT <= (A AND B) OR (A AND CIN) OR (B AND CIN); 
END SOMADOR_ARCH;