LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SOMADORPALAVRAS IS
PORT (
A,B : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
S : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
);
END SOMADORPALAVRAS;

ARCHITECTURE SUM OF SOMADORPALAVRAS IS

COMPONENT SOMADORCOMP IS
PORT (
A, B, CIN : IN STD_LOGIC;
S, COUT : OUT STD_LOGIC

);
END COMPONENT;

SIGNAL CARRY : STD_LOGIC_VECTOR(4 DOWNTO 0);

BEGIN

CARRY(0) <= '0';

SOMADOR1: SOMADORCOMP PORT MAP(
A => A(0),
B => B(0),
CIN => CARRY(0),
S => S(0),
COUT => CARRY(1)
);

SOMADOR2: SOMADORCOMP PORT MAP(
A => A(1),
B => B(1),
CIN => CARRY(1),
S => S(1),
COUT => CARRY(2)
);

SOMADOR3: SOMADORCOMP PORT MAP(
A => A(2),
B => B(2),
CIN => CARRY(2),
S => S(2),
COUT => CARRY(3)
);

SOMADOR4: SOMADORCOMP PORT MAP(
A => A(3),
B => B(3),
CIN => CARRY(3),
S => S(3),
COUT => CARRY(4)
);


S(4) <= CARRY(4);

END SUM;
