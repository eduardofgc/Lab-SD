LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY CONTADOR_100 IS
	PORT(CLK, RESET, ENABLE, LOAD: IN STD_LOGIC;
	     D_UN: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
	     D_DEZ: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
	     Q_UN: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
	     Q_DEZ: OUT STD_LOGIC_VECTOR (3 DOWNTO 0));
END CONTADOR_100;

ARCHITECTURE CONTADOR_100_ARCH OF CONTADOR_100 IS

COMPONENT CONTADOR10 IS
	PORT(CLK, RESET, ENABLE, RCI, LOAD: IN STD_LOGIC;
	     D: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
	     Q: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
	     RCO: OUT STD_LOGIC);
END COMPONENT;

SIGNAL UN_OUT: STD_LOGIC_VECTOR (3 DOWNTO 0);
SIGNAL DEZ_OUT: STD_LOGIC_VECTOR (3 DOWNTO 0);
SIGNAL CARRY: STD_LOGIC;

BEGIN

	UNIDADE: CONTADOR10 PORT MAP(CLK, RESET, ENABLE, '0', LOAD, D_UN, UN_OUT, CARRY);
	DEZENA: CONTADOR10 PORT MAP(CLK, RESET, CARRY, '0', LOAD, D_DEZ, DEZ_OUT, OPEN);

	Q_UN <= UN_OUT;
	Q_DEZ <= DEZ_OUT;

END CONTADOR_100_ARCH;
