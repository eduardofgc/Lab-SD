LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY TBSOMADOR IS
END ENTITY TBSOMADOR;

ARCHITECTURE TESTBENCH OF TBSOMADOR IS

COMPONENT GOLDENSOMADOR IS
PORT (
A, B : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
S : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
);
END COMPONENT;


SIGNAL A, B : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL S : STD_LOGIC_VECTOR(4 DOWNTO 0);

BEGIN

DUT: GOLDENSOMADOR PORT MAP (
A => A,
B => B,
S => S
);

ESTIMULOS: PROCESS
VARIABLE I : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
BEGIN
FOR count IN 0 TO 255 LOOP
A <= I(3 DOWNTO 0);
B <= I(7 DOWNTO 4);
WAIT FOR 500 NS;
I := STD_LOGIC_VECTOR(UNSIGNED(I) + 1);
END LOOP;


END PROCESS ESTIMULOS;

END ARCHITECTURE TESTBENCH;
