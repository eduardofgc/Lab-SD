LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY SOMADOR_ARITMETICO IS
	PORT(A: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
	     B: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
	     S: OUT STD_LOGIC_VECTOR (4 DOWNTO 0));
END ENTITY SOMADOR_ARITMETICO;

ARCHITECTURE SOMADOR_ARITMETICO_ARCH OF SOMADOR_ARITMETICO IS
BEGIN
	S <= ('0' & UNSIGNED(A)) + ('0' & UNSIGNED(B));
END ARCHITECTURE SOMADOR_ARITMETICO_ARCH;