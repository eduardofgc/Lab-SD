LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SOMADOR_COMPLETO IS
	PORT(A, B, CIN: IN STD_LOGIC;
	     S, COUT: OUT STD_LOGIC);
END ENTITY SOMADOR_COMPLETO;

ARCHITECTURE SOMADOR_COMPLETO_ARCH OF SOMADOR_COMPLETO IS
BEGIN
	S <= A XOR B XOR CIN;
	COUT <= (A AND B) OR (A AND CIN) OR (B AND CIN);
END ARCHITECTURE SOMADOR_COMPLETO_ARCH;
