LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MY_CIRCUIT3 IS
	PORT(A, B, C, D, E, F, G: IN STD_LOGIC;
	     Z: OUT STD_LOGIC);
END MY_CIRCUIT3;

ARCHITECTURE MY_CIRCUIT3_ARCH OF MY_CIRCUIT3 IS

	COMPONENT DECOD IS
		PORT (A: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		      B: OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
	END COMPONENT DECOD;

	COMPONENT MUX IS
		PORT (D: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		      S: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		      Y: OUT STD_LOGIC);
	END COMPONENT MUX;

	SIGNAL A1: STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL B1: STD_LOGIC_VECTOR (15 DOWNTO 0);

	SIGNAL D1: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL S1: STD_LOGIC_VECTOR (2 DOWNTO 0);
	SIGNAL Y1: STD_LOGIC;

BEGIN
	DEC_INST: DECOD PORT MAP(A => A1, B => B1);
	MUX_INST: MUX PORT MAP(D => D1, S => S1, Y => Y1);

	A1 <= A & B & C & D;
	D1 <= '1' & (B1(10) OR B1(11)) & '0' & (B1(9) OR B1(15)) & '1' & B1(7) & (B1(0) OR B1(15)) & '0';
	S1 <= E & F & G;
	Z <= Y1;

END MY_CIRCUIT3_ARCH;