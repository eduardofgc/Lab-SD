LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY CONTADOR10 IS
	PORT (CLK, RESET, ENABLE, RCI, LOAD: IN STD_LOGIC;
	      D: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	      Q: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
              RCO: OUT STD_LOGIC);
END CONTADOR10;

ARCHITECTURE CONTADOR_ARCH OF CONTADOR10 IS

	TYPE STATE IS(S0, S1, S2, S3, S4, S5, S6, S7, S8, S9);
	SIGNAL ESTADO_ATUAL, PROX_ESTADO, LOAD_ESTADO: STATE;

BEGIN

WITH D SELECT
	LOAD_ESTADO <= S0 WHEN "0000",
		       S1 WHEN "0001",
		       S2 WHEN "0010",
                       S3 WHEN "0011",
		       S4 WHEN "0100",
		       S5 WHEN "0101",
		       S6 WHEN "0110",
		       S7 WHEN "0111",
		       S8 WHEN "1000",
		       S9 WHEN "1001",
		       S0 WHEN OTHERS;

PROCESSO_SINCRONO: PROCESS(CLK)
BEGIN

IF RISING_EDGE(CLK) THEN
	ESTADO_ATUAL <= PROX_ESTADO;
END IF;

END PROCESS;

PROCESSO_COMBINACIONAL: PROCESS(ESTADO_ATUAL, RESET, ENABLE, RCI, LOAD, LOAD_ESTADO)
BEGIN

CASE ESTADO_ATUAL IS

	WHEN S0 =>
		Q <= "0000";
		RCO <= '1';
		
		IF (RESET = '1') THEN PROX_ESTADO <= S0;
		ELSIF (LOAD = '1') THEN PROX_ESTADO <= LOAD_ESTADO;
		ELSIF ((ENABLE = '0') AND (RCI = '0')) THEN PROX_ESTADO <= S1;
		ELSE PROX_ESTADO <= S0;
		END IF;

	WHEN S1 =>
		Q <= "0001";
		RCO <= '1';

		IF (RESET = '1') THEN PROX_ESTADO <= S0;
		ELSIF (LOAD = '1') THEN PROX_ESTADO <= LOAD_ESTADO;
		ELSIF ((ENABLE = '0') AND (RCI = '0')) THEN PROX_ESTADO <= S2;
		ELSE PROX_ESTADO <= S1;
		END IF;

	WHEN S2 =>
		Q <= "0010";
		RCO <= '1';

		IF (RESET = '1') THEN PROX_ESTADO <= S0;
		ELSIF (LOAD = '1') THEN PROX_ESTADO <= LOAD_ESTADO;
		ELSIF ((ENABLE = '0') AND (RCI = '0')) THEN PROX_ESTADO <= S3;
		ELSE PROX_ESTADO <= S2;
		END IF;

	WHEN S3 =>
		Q <= "0011";
		RCO <= '1';

		IF (RESET = '1') THEN PROX_ESTADO <= S0;
		ELSIF (LOAD = '1') THEN PROX_ESTADO <= LOAD_ESTADO;
		ELSIF ((ENABLE = '0') AND (RCI = '0')) THEN PROX_ESTADO <= S4;
		ELSE PROX_ESTADO <= S3;
		END IF;

	WHEN S4 =>
		Q <= "0100";
		RCO <= '1';

		IF (RESET = '1') THEN PROX_ESTADO <= S0;
		ELSIF (LOAD = '1') THEN PROX_ESTADO <= LOAD_ESTADO;
		ELSIF ((ENABLE = '0') AND (RCI = '0')) THEN PROX_ESTADO <= S5;
		ELSE PROX_ESTADO <= S4;
		END IF;

	WHEN S5 =>
		Q <= "0101";
		RCO <= '1';

		IF (RESET = '1') THEN PROX_ESTADO <= S0;
		ELSIF (LOAD = '1') THEN PROX_ESTADO <= LOAD_ESTADO;
		ELSIF ((ENABLE = '0') AND (RCI = '0')) THEN PROX_ESTADO <= S6;
		ELSE PROX_ESTADO <= S5;
		END IF;

	WHEN S6 =>
		Q <= "0110";
		RCO <= '1';

		IF (RESET = '1') THEN PROX_ESTADO <= S0;
		ELSIF (LOAD = '1') THEN PROX_ESTADO <= LOAD_ESTADO;
		ELSIF ((ENABLE = '0') AND (RCI = '0')) THEN PROX_ESTADO <= S7;
		ELSE PROX_ESTADO <= S6;
		END IF;

	WHEN S7 =>
		Q <= "0111";
		RCO <= '1';

		IF (RESET = '1') THEN PROX_ESTADO <= S0;
		ELSIF (LOAD = '1') THEN PROX_ESTADO <= LOAD_ESTADO;
		ELSIF ((ENABLE = '0') AND (RCI = '0')) THEN PROX_ESTADO <= S8;
		ELSE PROX_ESTADO <= S7;
		END IF;

	WHEN S8 =>
		Q <= "1000";
		RCO <= '1';

		IF (RESET = '1') THEN PROX_ESTADO <= S0;
		ELSIF (LOAD = '1') THEN PROX_ESTADO <= LOAD_ESTADO;
		ELSIF ((ENABLE = '0') AND (RCI = '0')) THEN PROX_ESTADO <= S9;
		ELSE PROX_ESTADO <= S8;
		END IF;

	WHEN S9 =>
		Q <= "1001";
		RCO <= '0';

		IF (RESET = '1') THEN PROX_ESTADO <= S0;
		ELSIF (LOAD = '1') THEN PROX_ESTADO <= LOAD_ESTADO;
		ELSIF ((ENABLE = '0') AND (RCI = '0')) THEN PROX_ESTADO <= S0;
		ELSE PROX_ESTADO <= S9;
		END IF;

	WHEN OTHERS =>
		Q <= "0000";
		RCO <= '1';

		IF (RESET = '1') THEN PROX_ESTADO <= S0;
		ELSIF (LOAD = '1') THEN PROX_ESTADO <= LOAD_ESTADO;
		ELSIF ((ENABLE = '0') AND (RCI = '0')) THEN PROX_ESTADO <= S1;
		ELSE PROX_ESTADO <= S0;
		END IF;
END CASE;
END PROCESS;

END CONTADOR_ARCH;
