LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY TESTBENCH_SOMADOR IS
END ENTITY TESTBENCH_SOMADOR;

ARCHITECTURE TESTBENCH_SOMADOR_ARCH OF TESTBENCH_SOMADOR IS

COMPONENT TB_SOMADOR_4BITS IS
	PORT(A: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
	     B: OUT STD_LOGIC_VECTOR (3 DOWNTO 0));
END COMPONENT TB_SOMADOR_4BITS;

COMPONENT SOMADOR_PALAVRAS_4BITS IS
	PORT(A: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
	     B: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
	     S: OUT STD_LOGIC_VECTOR (4 DOWNTO 0));
END COMPONENT SOMADOR_PALAVRAS_4BITS;

COMPONENT SOMADOR_ARITMETICO IS
	PORT(A: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
	     B: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
	     S: OUT STD_LOGIC_VECTOR (4 DOWNTO 0));
END COMPONENT SOMADOR_ARITMETICO;

SIGNAL A_TESTBENCH, B_TESTBENCH: STD_LOGIC_VECTOR (3 DOWNTO 0);
SIGNAL S_TESTBENCH, S_TESTBENCH_ARITMETICO: STD_LOGIC_VECTOR (4 DOWNTO 0);

BEGIN

	TESTBENCH: COMPONENT TB_SOMADOR_4BITS
		PORT MAP(A => A_TESTBENCH, B => B_TESTBENCH);

	EX_SOMADOR_PALAVRAS_4BITS: COMPONENT SOMADOR_PALAVRAS_4BITS
		PORT MAP(A => A_TESTBENCH, B => B_TESTBENCH, S => S_TESTBENCH);

	EX_SOMADOR_ARITMETICO: COMPONENT SOMADOR_ARITMETICO
		PORT MAP(A => A_TESTBENCH, B => B_TESTBENCH, S => S_TESTBENCH_ARITMETICO);

	PROCESSO_COMPARACIONAL: PROCESS(A_TESTBENCH, B_TESTBENCH)
	BEGIN
		IF S_TESTBENCH /= S_TESTBENCH_ARITMETICO THEN
			REPORT "INCONSISTENCIA. S_TESTBENCH = " & INTEGER'IMAGE(to_integer(unsigned(S_TESTBENCH))) & " E S_TESTBENCH_ARITMETICO = " & INTEGER'IMAGE(to_integer(unsigned(S_TESTBENCH_ARITMETICO)));
		END IF;
	END PROCESS;

END ARCHITECTURE TESTBENCH_SOMADOR_ARCH;
	
