LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE STD.TEXTIO.ALL;
USE IEEE.NUMERIC_STD;

ENTITY MAQUINA_DE_ESTADOS IS
	PORT(A: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
	     CLOCK, RESET: IN STD_LOGIC;
	     P, T25, T50: OUT STD_LOGIC);
END MAQUINA_DE_ESTADOS;

ARCHITECTURE MAQUINA_DE_ESTADOS_ARCH OF MAQUINA_DE_ESTADOS IS

TYPE ESTADOS IS (INIT, S25, S50, S75, S100, S125, D25, D50, D75);

SIGNAL ESTADO_ATUAL, PROX_ESTADO : ESTADOS;

BEGIN

	PROCESSO : PROCESS(CLOCK, RESET)
	BEGIN

	IF (RESET = '1') THEN
		ESTADO_ATUAL <= INIT;
	ELSIF (RISING_EDGE(CLOCK)) THEN
		ESTADO_ATUAL <= PROX_ESTADO;
	END IF;

END PROCESS PROCESSO;

PROCESSO_COMB : PROCESS(ESTADO_ATUAL, A)
BEGIN

CASE ESTADO_ATUAL IS

WHEN INIT => P <= '0'; T25 <= '0'; T50 <= '0';

IF A = "00" THEN PROX_ESTADO <= INIT;
ELSIF A = "01" THEN PROX_ESTADO <= S25;
ELSIF A = "10" THEN PROX_ESTADO <= S50;
ELSIF A = "11" THEN PROX_ESTADO <= INIT;

END IF;

WHEN S25 => P <= '0'; T25 <= '0'; T50 <= '0';

IF A = "00" THEN PROX_ESTADO <= S25;
ELSIF A = "01" THEN PROX_ESTADO <= S50;
ELSIF A = "10" THEN PROX_ESTADO <= S75;
ELSIF A = "11" THEN PROX_ESTADO <= D25;

END IF;

WHEN S50 => P <= '0'; T25 <= '0'; T50 <= '0';

IF A = "00" THEN PROX_ESTADO <= S50;
ELSIF A = "01" THEN PROX_ESTADO <= S75;
ELSIF A = "10" THEN PROX_ESTADO <= S100;
ELSIF A = "11" THEN PROX_ESTADO <= D50;

END IF;

WHEN S75 => P <= '0'; T25 <= '0'; T50 <= '0';

IF A = "00" THEN PROX_ESTADO <= S75;
ELSIF A = "01" THEN PROX_ESTADO <= S100;
ELSIF A = "10" THEN PROX_ESTADO <= S125;
ELSIF A = "11" THEN PROX_ESTADO <= D75;

END IF;

WHEN S100 => P <= '1'; T25 <= '0'; T50 <= '0';

IF A = "00" THEN PROX_ESTADO <= INIT;
ELSIF A = "01" THEN PROX_ESTADO <= INIT;
ELSIF A = "10" THEN PROX_ESTADO <= INIT;
ELSIF A = "11" THEN PROX_ESTADO <= INIT;

END IF;

WHEN S125 => P <= '1'; T25 <= '1'; T50 <= '0';

IF A = "00" THEN PROX_ESTADO <= INIT;
ELSIF A = "01" THEN PROX_ESTADO <= INIT;
ELSIF A = "10" THEN PROX_ESTADO <= INIT;
ELSIF A = "11" THEN PROX_ESTADO <= INIT;

END IF;

WHEN D25 => P <= '0'; T25 <= '1'; T50 <= '0';

IF A = "00" THEN PROX_ESTADO <= INIT;
ELSIF A = "01" THEN PROX_ESTADO <= S25;
ELSIF A = "10" THEN PROX_ESTADO <= S50;
ELSIF A = "11" THEN PROX_ESTADO <= INIT;

END IF;

WHEN D50 => P <= '0'; T25 <= '0'; T50 <= '1';

IF A = "00" THEN PROX_ESTADO <= INIT;
ELSIF A = "01" THEN PROX_ESTADO <= S25;
ELSIF A = "10" THEN PROX_ESTADO <= S50;
ELSIF A = "11" THEN PROX_ESTADO <= INIT;

END IF;

WHEN D75 => P <= '0'; T25 <= '1'; T50 <= '1';

IF A = "00" THEN PROX_ESTADO <= INIT;
ELSIF A = "01" THEN PROX_ESTADO <= S25;
ELSIF A = "10" THEN PROX_ESTADO <= S50;
ELSIF A = "11" THEN PROX_ESTADO <= INIT;

END IF;

END CASE;

END PROCESS PROCESSO_COMB;

END MAQUINA_DE_ESTADOS_ARCH;